module sub1 #(
	parameter DATA_WIDTH = 1'b0
)(
	input  clk,
	input  rst,
	output  intr);

	//Wire define for this module.

	//Wire define for sub module.

	//Wire sub module connect to this module and inter module connect.

	//Wire this module connect to sub module.

	//module inst.

endmodule