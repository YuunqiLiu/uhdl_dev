module sub1 (
	input  clk,
	input  rst,
	output  intr);

	//Wire define for this module.

	//Wire define for sub module.

	//Wire sub module connect to this module and inter module connect.
	assign sub1_clk = clk;

	//Wire this module connect to sub module.

	//module inst.

endmodule