module AXICrossbar(
    input  acr_clk,
    input  acr_rst,
    input [31:0] axii0_awaddr,
    input [3:0] axii0_awlen,
    input [2:0] axii0_awsize,
    input [1:0] axii0_awburst,
    input  axii0_awlock,
    input [3:0] axii0_awcache,
    input [2:0] axii0_awprot,
    input  axii0_awvalid,
    output  axii0_awready,
    input [63:0] axii0_wdata,
    input [7:0] axii0_wstrb,
    input  axii0_wlast,
    input  axii0_wvalid,
    output  axii0_wready,
    output [7:0] axii0_bid,
    output [1:0] axii0_bresp,
    output  axii0_bvalid,
    input  axii0_bready,
    input [7:0] axii0_arid,
    input [31:0] axii0_araddr,
    input [3:0] axii0_arlen,
    input [2:0] axii0_arsize,
    input [1:0] axii0_arburst,
    input  axii0_arlock,
    input [3:0] axii0_arcache,
    input [2:0] axii0_arprot,
    input  axii0_arvalid,
    output  axii0_arready,
    output [7:0] axii0_rid,
    output [63:0] axii0_rdata,
    output [1:0] axii0_rresp,
    output  axii0_rlast,
    output  axii0_rvalid,
    input  axii0_rready,
    input [31:0] axii1_awaddr,
    input [3:0] axii1_awlen,
    input [2:0] axii1_awsize,
    input [1:0] axii1_awburst,
    input  axii1_awlock,
    input [3:0] axii1_awcache,
    input [2:0] axii1_awprot,
    input  axii1_awvalid,
    output  axii1_awready,
    input [63:0] axii1_wdata,
    input [7:0] axii1_wstrb,
    input  axii1_wlast,
    input  axii1_wvalid,
    output  axii1_wready,
    output [7:0] axii1_bid,
    output [1:0] axii1_bresp,
    output  axii1_bvalid,
    input  axii1_bready,
    input [7:0] axii1_arid,
    input [31:0] axii1_araddr,
    input [3:0] axii1_arlen,
    input [2:0] axii1_arsize,
    input [1:0] axii1_arburst,
    input  axii1_arlock,
    input [3:0] axii1_arcache,
    input [2:0] axii1_arprot,
    input  axii1_arvalid,
    output  axii1_arready,
    output [7:0] axii1_rid,
    output [63:0] axii1_rdata,
    output [1:0] axii1_rresp,
    output  axii1_rlast,
    output  axii1_rvalid,
    input  axii1_rready,
    input [31:0] axii2_awaddr,
    input [3:0] axii2_awlen,
    input [2:0] axii2_awsize,
    input [1:0] axii2_awburst,
    input  axii2_awlock,
    input [3:0] axii2_awcache,
    input [2:0] axii2_awprot,
    input  axii2_awvalid,
    output  axii2_awready,
    input [63:0] axii2_wdata,
    input [7:0] axii2_wstrb,
    input  axii2_wlast,
    input  axii2_wvalid,
    output  axii2_wready,
    output [7:0] axii2_bid,
    output [1:0] axii2_bresp,
    output  axii2_bvalid,
    input  axii2_bready,
    input [7:0] axii2_arid,
    input [31:0] axii2_araddr,
    input [3:0] axii2_arlen,
    input [2:0] axii2_arsize,
    input [1:0] axii2_arburst,
    input  axii2_arlock,
    input [3:0] axii2_arcache,
    input [2:0] axii2_arprot,
    input  axii2_arvalid,
    output  axii2_arready,
    output [7:0] axii2_rid,
    output [63:0] axii2_rdata,
    output [1:0] axii2_rresp,
    output  axii2_rlast,
    output  axii2_rvalid,
    input  axii2_rready,
    input [31:0] axii3_awaddr,
    input [3:0] axii3_awlen,
    input [2:0] axii3_awsize,
    input [1:0] axii3_awburst,
    input  axii3_awlock,
    input [3:0] axii3_awcache,
    input [2:0] axii3_awprot,
    input  axii3_awvalid,
    output  axii3_awready,
    input [63:0] axii3_wdata,
    input [7:0] axii3_wstrb,
    input  axii3_wlast,
    input  axii3_wvalid,
    output  axii3_wready,
    output [7:0] axii3_bid,
    output [1:0] axii3_bresp,
    output  axii3_bvalid,
    input  axii3_bready,
    input [7:0] axii3_arid,
    input [31:0] axii3_araddr,
    input [3:0] axii3_arlen,
    input [2:0] axii3_arsize,
    input [1:0] axii3_arburst,
    input  axii3_arlock,
    input [3:0] axii3_arcache,
    input [2:0] axii3_arprot,
    input  axii3_arvalid,
    output  axii3_arready,
    output [7:0] axii3_rid,
    output [63:0] axii3_rdata,
    output [1:0] axii3_rresp,
    output  axii3_rlast,
    output  axii3_rvalid,
    input  axii3_rready,
    input [31:0] axii4_awaddr,
    input [3:0] axii4_awlen,
    input [2:0] axii4_awsize,
    input [1:0] axii4_awburst,
    input  axii4_awlock,
    input [3:0] axii4_awcache,
    input [2:0] axii4_awprot,
    input  axii4_awvalid,
    output  axii4_awready,
    input [63:0] axii4_wdata,
    input [7:0] axii4_wstrb,
    input  axii4_wlast,
    input  axii4_wvalid,
    output  axii4_wready,
    output [7:0] axii4_bid,
    output [1:0] axii4_bresp,
    output  axii4_bvalid,
    input  axii4_bready,
    input [7:0] axii4_arid,
    input [31:0] axii4_araddr,
    input [3:0] axii4_arlen,
    input [2:0] axii4_arsize,
    input [1:0] axii4_arburst,
    input  axii4_arlock,
    input [3:0] axii4_arcache,
    input [2:0] axii4_arprot,
    input  axii4_arvalid,
    output  axii4_arready,
    output [7:0] axii4_rid,
    output [63:0] axii4_rdata,
    output [1:0] axii4_rresp,
    output  axii4_rlast,
    output  axii4_rvalid,
    input  axii4_rready,
    output [31:0] axio0_awaddr,
    output [3:0] axio0_awlen,
    output [2:0] axio0_awsize,
    output [1:0] axio0_awburst,
    output  axio0_awlock,
    output [3:0] axio0_awcache,
    output [2:0] axio0_awprot,
    output  axio0_awvalid,
    input  axio0_awready,
    output [63:0] axio0_wdata,
    output [7:0] axio0_wstrb,
    output  axio0_wlast,
    output  axio0_wvalid,
    input  axio0_wready,
    input [7:0] axio0_bid,
    input [1:0] axio0_bresp,
    input  axio0_bvalid,
    output  axio0_bready,
    output [7:0] axio0_arid,
    output [31:0] axio0_araddr,
    output [3:0] axio0_arlen,
    output [2:0] axio0_arsize,
    output [1:0] axio0_arburst,
    output  axio0_arlock,
    output [3:0] axio0_arcache,
    output [2:0] axio0_arprot,
    output  axio0_arvalid,
    input  axio0_arready,
    input [7:0] axio0_rid,
    input [63:0] axio0_rdata,
    input [1:0] axio0_rresp,
    input  axio0_rlast,
    input  axio0_rvalid,
    output  axio0_rready,
    output [31:0] axio1_awaddr,
    output [3:0] axio1_awlen,
    output [2:0] axio1_awsize,
    output [1:0] axio1_awburst,
    output  axio1_awlock,
    output [3:0] axio1_awcache,
    output [2:0] axio1_awprot,
    output  axio1_awvalid,
    input  axio1_awready,
    output [63:0] axio1_wdata,
    output [7:0] axio1_wstrb,
    output  axio1_wlast,
    output  axio1_wvalid,
    input  axio1_wready,
    input [7:0] axio1_bid,
    input [1:0] axio1_bresp,
    input  axio1_bvalid,
    output  axio1_bready,
    output [7:0] axio1_arid,
    output [31:0] axio1_araddr,
    output [3:0] axio1_arlen,
    output [2:0] axio1_arsize,
    output [1:0] axio1_arburst,
    output  axio1_arlock,
    output [3:0] axio1_arcache,
    output [2:0] axio1_arprot,
    output  axio1_arvalid,
    input  axio1_arready,
    input [7:0] axio1_rid,
    input [63:0] axio1_rdata,
    input [1:0] axio1_rresp,
    input  axio1_rlast,
    input  axio1_rvalid,
    output  axio1_rready,
    output [31:0] axio2_awaddr,
    output [3:0] axio2_awlen,
    output [2:0] axio2_awsize,
    output [1:0] axio2_awburst,
    output  axio2_awlock,
    output [3:0] axio2_awcache,
    output [2:0] axio2_awprot,
    output  axio2_awvalid,
    input  axio2_awready,
    output [63:0] axio2_wdata,
    output [7:0] axio2_wstrb,
    output  axio2_wlast,
    output  axio2_wvalid,
    input  axio2_wready,
    input [7:0] axio2_bid,
    input [1:0] axio2_bresp,
    input  axio2_bvalid,
    output  axio2_bready,
    output [7:0] axio2_arid,
    output [31:0] axio2_araddr,
    output [3:0] axio2_arlen,
    output [2:0] axio2_arsize,
    output [1:0] axio2_arburst,
    output  axio2_arlock,
    output [3:0] axio2_arcache,
    output [2:0] axio2_arprot,
    output  axio2_arvalid,
    input  axio2_arready,
    input [7:0] axio2_rid,
    input [63:0] axio2_rdata,
    input [1:0] axio2_rresp,
    input  axio2_rlast,
    input  axio2_rvalid,
    output  axio2_rready
);



endmodule