module Adder (
	input        in1,
	input        in2,
	output [1:0] out);

	//Wire define for this module.

	//Wire define for sub module.

	//Wire sub module connect to this module and inter module connect.
	assign out = (in1 + in2);
	

	//Wire this module connect to sub module.

	//module inst.

endmodule