module clk_divider_1600_to_150 (
	input  clk_in,
	output  clk_out);

	//Wire define for this module.

	//Wire define for sub module.

	//Wire sub module connect to this module and inter module connect.

	//Wire this module connect to sub module.

	//module inst.

endmodule