module AISRAM(
    input  acr_clk,
    input  acr_rst,
    input [31:0] axi_awaddr,
    input [3:0] axi_awlen,
    input [2:0] axi_awsize,
    input [1:0] axi_awburst,
    input  axi_awlock,
    input [3:0] axi_awcache,
    input [2:0] axi_awprot,
    input  axi_awvalid,
    output  axi_awready,
    input [63:0] axi_wdata,
    input [7:0] axi_wstrb,
    input  axi_wlast,
    input  axi_wvalid,
    output  axi_wready,
    output [7:0] axi_bid,
    output [1:0] axi_bresp,
    output  axi_bvalid,
    input  axi_bready,
    input [7:0] axi_arid,
    input [31:0] axi_araddr,
    input [3:0] axi_arlen,
    input [2:0] axi_arsize,
    input [1:0] axi_arburst,
    input  axi_arlock,
    input [3:0] axi_arcache,
    input [2:0] axi_arprot,
    input  axi_arvalid,
    output  axi_arready,
    output [7:0] axi_rid,
    output [63:0] axi_rdata,
    output [1:0] axi_rresp,
    output  axi_rlast,
    output  axi_rvalid,
    input  axi_rready
);



endmodule